module rotating_mode_cordic(
    input [11:0]x_value,
    input [11:0]y_value,
    input [6:0]angle, // [6]Signed 1-bit, [5:0]Data 6-bit  +99 ~ -99
    output [11:0]x_out,
    output [11:0]y_out
);

// iteration = 8



endmodule