module local_oscillator_nsin(
    input clk_8megahz,
    input rst_n,
    input wire signed [13:0] filtered_data,
    output reg signed [13:0] lo_nsin_data
);

endmodule