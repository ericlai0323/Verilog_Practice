module map(mode, pattern, map1, map2, map3, map4, map5, map6, map7, map8);

output reg [7:0]map1, map2, map3, map4, map5, map6, map7, map8;
input [2:0]pattern; 
input [1:0]mode;

always@(mode or pattern)
begin
    case(mode)
    2'd0:
    begin
        case(pattern)
            //walk
            4'd0:
            begin 
                map1 <= 8'b0011_1000;
                map2 <= 8'b0011_0000;
                map3 <= 8'b0001_1110;
                map4 <= 8'b0011_1001;
                map5 <= 8'b0100_1000;
                map6 <= 8'b0001_0100;
                map7 <= 8'b0010_0010; 
                map8 <= 8'b0110_0001;
            end
            4'd1:
            begin 
                map1 <= 8'b0011_1000;
                map2 <= 8'b0011_0000;
                map3 <= 8'b0001_1110;
                map4 <= 8'b0011_1011;
                map5 <= 8'b0110_1000;
                map6 <= 8'b0001_0100;
                map7 <= 8'b0010_0100; 
                map8 <= 8'b0010_0010;
            end
            4'd2:
            begin 
                map1 <= 8'b0011_1000;
                map2 <= 8'b0011_0000;
                map3 <= 8'b0001_1100;
                map4 <= 8'b0001_1010;
                map5 <= 8'b0010_1010;
                map6 <= 8'b0001_0100;
                map7 <= 8'b0010_0100; 
                map8 <= 8'b0010_0010;
            end
            4'd3:
            begin 
                map1 <= 8'b0011_1000;
                map2 <= 8'b0011_0000;
                map3 <= 8'b0001_1000;
                map4 <= 8'b0001_1100;
                map5 <= 8'b0001_1000;
                map6 <= 8'b0000_1100;
                map7 <= 8'b0001_0100; 
                map8 <= 8'b0010_0100;
            end
            4'd4:
            begin 
                map1 <= 8'b0011_1000;
                map2 <= 8'b0011_0000;
                map3 <= 8'b0001_1000;
                map4 <= 8'b0001_1000;
                map5 <= 8'b0001_1000;
                map6 <= 8'b0000_1100;
                map7 <= 8'b0000_1100; 
                map8 <= 8'b0000_0100;
            end
            4'd5:
            begin 
                map1 <= 8'b0011_1000;
                map2 <= 8'b0011_0000;
                map3 <= 8'b0001_1100;
                map4 <= 8'b0001_1000;
                map5 <= 8'b0011_1000;
                map6 <= 8'b0000_1100;
                map7 <= 8'b0001_0100; 
                map8 <= 8'b0001_0010;
            end
            4'd6:
            begin 
                map1 <= 8'b0011_1000;
                map2 <= 8'b0011_0000;
                map3 <= 8'b0001_1100;
                map4 <= 8'b0011_1010;
                map5 <= 8'b0101_1000;
                map6 <= 8'b0000_1000;
                map7 <= 8'b0001_0100; 
                map8 <= 8'b0010_0010;
            end
            4'd7:
            begin 
                map1 <= 8'b0011_1000;
                map2 <= 8'b0011_0000;
                map3 <= 8'b0001_1110;
                map4 <= 8'b0111_1001;
                map5 <= 8'b1001_1000;
                map6 <= 8'b0001_1000;
                map7 <= 8'b0010_0100; 
                map8 <= 8'b0100_0010;
            end
        endcase
    end
    //run
    2'd1:
    begin
        case(pattern)
            4'd0:
            begin 
                map1 <= 8'b0110_0000;	                map2 <= 8'b0110_0000;
                map3 <= 8'b0011_0000;
                map4 <= 8'b0111_1000;
                map5 <= 8'b0001_1000;
                map6 <= 8'b0011_0100;
                map7 <= 8'b0010_0010; 
                map8 <= 8'b0110_0110;
            end
            4'd1:
            begin 
                map1 <= 8'b0110_0000;
                map2 <= 8'b0110_0000;
                map3 <= 8'b0011_0000;
                map4 <= 8'b0111_1100;
                map5 <= 8'b0101_1010;
                map6 <= 8'b0011_0100;
                map7 <= 8'b0110_0010; 
                map8 <= 8'b0100_0010;
            end
            4'd2:
            begin 
                map1 <= 8'b0110_0000;
                map2 <= 8'b0110_0000;
                map3 <= 8'b0011_0000;
                map4 <= 8'b0111_1100;
                map5 <= 8'b1011_0010;
                map6 <= 8'b0001_1000;
                map7 <= 8'b0110_0110; 
                map8 <= 8'b0000_0010;
            end
            4'd3:
            begin 
                map1 <= 8'b1100_0000;
                map2 <= 8'b1100_0000;
                map3 <= 8'b0111_1000;
                map4 <= 8'b0110_0100;
                map5 <= 8'b1011_0000;
                map6 <= 8'b0010_1000;
                map7 <= 8'b1100_0110; 
                map8 <= 8'b0000_0010;
            end
            4'd4:
            begin 
                map1 <= 8'b1100_0000;
                map2 <= 8'b1100_0000;
                map3 <= 8'b0110_0000;
                map4 <= 8'b0111_1000;
                map5 <= 8'b1011_0100;
                map6 <= 8'b0011_1010;
                map7 <= 8'b0010_0110; 
                map8 <= 8'b1110_0010;
            end
            4'd5:
            begin 
                map1 <= 8'b1100_0000;
                map2 <= 8'b1100_0000;
                map3 <= 8'b0110_0000;
                map4 <= 8'b0111_1000;
                map5 <= 8'b1011_0100;
                map6 <= 8'b0011_0010;
                map7 <= 8'b0100_1100; 
                map8 <= 8'b1100_0100;
            end
            4'd6:
            begin 
                map1 <= 8'b1100_0000;
                map2 <= 8'b1100_0000;
                map3 <= 8'b0110_0000;
                map4 <= 8'b0111_1000;
                map5 <= 8'b0111_0100;
                map6 <= 8'b0011_0000;
                map7 <= 8'b0101_1000; 
                map8 <= 8'b0010_1000;
            end
            4'd7:
            begin 
                map1 <= 8'b0110_0000;
                map2 <= 8'b0110_0000;
                map3 <= 8'b0011_0000;
                map4 <= 8'b0011_1000;
                map5 <= 8'b0001_1000;
                map6 <= 8'b0001_0100;
                map7 <= 8'b0001_1100; 
                map8 <= 8'b0000_0100;
            end
        endcase
    end
    //stop
    2'd2:
    begin
        case(pattern)
            4'd0:
            begin 
                map1 <= 8'b0001_1000;
                map2 <= 8'b0001_1000;
                map3 <= 8'b0011_1100;
                map4 <= 8'b0101_1010;
                map5 <= 8'b0101_1010;
                map6 <= 8'b0001_1000;
                map7 <= 8'b0010_0100; 
                map8 <= 8'b0110_0110;
            end
        endcase
    end
    endcase
end

endmodule

