library verilog;
use verilog.vl_types.all;
entity top_bcd is
    port(
        clk_50megahz    : in     vl_logic;
        sw_a            : in     vl_logic_vector(3 downto 0);
        sw_b            : in     vl_logic_vector(3 downto 0);
        sw_mode         : in     vl_logic_vector(1 downto 0);
        flag_n          : in     vl_logic;
        rst_n           : in     vl_logic;
        sw_a_led        : out    vl_logic_vector(3 downto 0);
        sw_b_led        : out    vl_logic_vector(3 downto 0);
        sw_mode_led     : out    vl_logic_vector(1 downto 0);
        key_flag_n      : out    vl_logic;
        key_rst_n       : out    vl_logic;
        bcd_a_0_0       : out    vl_logic;
        bcd_a_0_1       : out    vl_logic;
        bcd_a_0_2       : out    vl_logic;
        bcd_a_0_3       : out    vl_logic;
        bcd_a_1_0       : out    vl_logic;
        bcd_a_1_1       : out    vl_logic;
        bcd_a_1_2       : out    vl_logic;
        bcd_a_1_3       : out    vl_logic;
        bcd_b_0_0       : out    vl_logic;
        bcd_b_0_1       : out    vl_logic;
        bcd_b_0_2       : out    vl_logic;
        bcd_b_0_3       : out    vl_logic;
        bcd_b_1_0       : out    vl_logic;
        bcd_b_1_1       : out    vl_logic;
        bcd_b_1_2       : out    vl_logic;
        bcd_b_1_3       : out    vl_logic;
        bcd_result_0_0  : out    vl_logic;
        bcd_result_0_1  : out    vl_logic;
        bcd_result_0_2  : out    vl_logic;
        bcd_result_0_3  : out    vl_logic;
        bcd_result_1_0  : out    vl_logic;
        bcd_result_1_1  : out    vl_logic;
        bcd_result_1_2  : out    vl_logic;
        bcd_result_1_3  : out    vl_logic;
        bcd_result_2_0  : out    vl_logic;
        bcd_result_2_1  : out    vl_logic;
        bcd_result_2_2  : out    vl_logic;
        bcd_result_2_3  : out    vl_logic;
        bcd_result_3_0  : out    vl_logic;
        bcd_result_3_1  : out    vl_logic;
        bcd_result_3_2  : out    vl_logic;
        bcd_result_3_3  : out    vl_logic
    );
end top_bcd;
